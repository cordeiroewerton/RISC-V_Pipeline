module Instr_Mem(input logic[7:0] A, output logic[31:0] RD);
	always_comb begin
		case(A)
			8'h00: RD = 32'b000000_00000_00000_00000_00000_000000;
			8'h04: RD = 32'b00000000011100000000000010010011;
			8'h08: RD = 32'b00000000001100000000000110010011;
			8'h0C: RD = 32'b11111111111100000000000100010011;
			8'h10: RD = 32'b00000000000100010000000100010011;
			8'h14: RD = 32'b00000000001100010010001110110011;
			8'h18: RD = 32'b11111110001000001000101011100011;
			8'h1C: RD = 32'b11111110000000000000101011100011;
			default: RD = 32'b000000_00000_00000_00000_00000_000000;
		endcase
	end
endmodule 
